module TestBench(FIFO_IF.TEST fifo_if);
    
endmodule