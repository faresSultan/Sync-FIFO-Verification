module tb(FIFO_IF.TEST fifo_if);
    
endmodule