package FIFO_coverage_pkg;

    class FIFO_coverage;

        
        
    endclass
endpackage